package defs;

	typedef enum logic [1:0]
	{
		ADD = 2'b00,
		SUB = 2'b01,
		AND = 2'b10,
		NOT = 2'b11
	} op_code_e;
	
endpackage
