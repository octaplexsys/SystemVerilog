module top (
	input		logic [ 2**N - 1 : 0 ]	line,
	output	logic [ N - 1 : 0 ]		code
	);
	
	
endmodule

module #(parameter WIDTH = 4) coder (
	input		logic [ 2**WIDTH - 1 : 0 ]	line,
	output	logic [ WIDTH - 1 : 0 ]		code
	);
	
	assign code
	
	
endmodule
