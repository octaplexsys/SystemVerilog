module UART_tx (
	input 	logic 				clk_i,
	input 	logic 				a_reset_i,
	input	logic				tx,
	input 	logic	[ 7 : 0 ]	tx_data,
	input	logic				tx_data_load_strobe
	);

endmodule // UART_tx
